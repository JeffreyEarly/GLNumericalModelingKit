netcdf tst_utf8 {
dimensions:
	Καλημέρα = 18 ;
variables:
	char Καλημέρα(Καλημέρα) ;
		Καλημέρα:units = "Καλημέρα" ;
data:

 Καλημέρα = "\316\232\316\261\316\273\316\267\316\274\341\275\263\317\201\316\261" ;
}
